library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;
    use ieee.std_logic_arith.all;

entity rom is
    port (
        ce      :in  std_logic;                      -- Chip Enable
        read_en :in  std_logic;                      -- Read Enable
        address :in  std_logic_vector (31 downto 0); -- Address input
        data    :out std_logic_vector (31 downto 0)  -- Data output
    );
end entity;
architecture rom_behavior of rom is

begin
--      func7     r2     r1     func3   rd      opcode
--mult 0000001  01011  01010    000   00101    0110011
  
--					         x5		REG Address
--       imm[11:5]     rs2        rs1       010   imm[4:0]      opcode
-- sw    0000000      00101      00010      010    00000     0100011

--       imm[11:5]     rs2        rs1       010   imm[4:0]      opcode
--																					0000011
       
    process (read_en, address) begin
        if (read_en = '1') then
            case (address) is
					--when x"00000000"   => data <= "00000000001000000000010100010011"; --addi x10 x0 2
               --when x"00000004"   => data <= "00000000101000000000010110010011"; --addi x11 x0 10 --li a1,10
               --when x"00000008"   => data <= "00000010101101010000001010110011"; --mult x5, x11 x10 --salva no x5
               --when x"0000000C"   => data <= "11111110101101010001111011100011"; --bne x10 x11 -4
               --when x"00000010"   => data <= "11111110101101010100100011100011"; --blt x10 x11 -16
               --when x"00000014"   => data <= "00000000101000000000010100010011"; --addi x10 x0 10
					-----------------------------------------------------------------------------------
					-----------------------------------------------------------------------------------
					--when x"00000000"   => data <= "00000000000000000000010100010011"; --addi x10 x0 0
               --when x"00000004"   => data <= "00000000101000000000010110010011"; --addi x11 x0 10 --li a1,10
               --when x"00000008"   => data <= "00000000000101010000010100010011"; --addi x10 x10 1
               --when x"0000000C"   => data <= "11111110101101010001111011100011"; --bne x10 x11 -4
               --when x"00000010"   => data <= "11111110101101010100100011100011"; --blt x10 x11 -16
					--when x"00000014"   => data <= "00000000001001110000011100010011"; --addi x14 x14 2
					--when x"00000018"   => data <= "11111110111001010001111011100011"; --bne x10 x14 -4
               --when x"00000014"   => data <= "00000000101000000000010100010011"; --addi x10 x0 10
					-----------------------------------------------------------------------------------
					-----------------------------------------------------------------------------------
					--when x"00000000"   => data <= "00000000000100000000010100010011";--addi x10 x0 1
               --when x"00000004"   => data <= "11111110010000010000000100010011";--addi x2 x2 -28
               --when x"00000008"   => data <= "00000000101000010010011000100011"; --sw x10 12(x2)
               --when x"0000000C"   => data <= "00000000110000010010011000000011"; --lw x12 12(x2)
               --when x"00000010"   => data <= "00000000110000010010011010000011"; --lw x13 12(x2)
					--when x"00000014"   => data <= "00000000101000000000010100010011"; --addi x10 x0 10
					-----------------------------------------------------------------------------------
					-----------------------------------------------------------------------------------
					when x"00000000"   => data <= "00000000000000000000000100010011"; --addi x2 x0 0
               when x"00000004"   => data <= "00000000010100000000001010010011"; --addi x5 x0 5
               when x"00000008"   => data <= "00000000010100010010000000100011"; --sw x5 0(x2)
               when x"0000000C"   => data <= "00000000000000010010010100000011"; --lw x10 0(x2)
               when x"00000010"   => data <= "00000000101000000000010110010011"; --addi x11 x0 10
               when x"00000014"   => data <= "00000000001000000000010100010011"; --addi x10 x0 2
					when x"00000018"   => data <= "00000010101101010000001010110011"; --mult x5, x11 x10
               when x"0000001C"   => data <= "11111110010000010000000100010011"; --addi x2 x2 -28
               when x"00000020"   => data <= "00000000101000010010011000100011"; --sw x10 12(x2)
               when x"00000024"   => data <= "00000000110000010010011000000011"; --lw x12 12(x2)
               when x"00000028"   => data <= "00000000000000000000010100010011"; --addi x10 x0 0
               when x"0000002C"   => data <= "00000000101000000000010110010011"; --addi x11 x0 10
               when x"00000030"   => data <= "00000000000101010000010100010011"; --addi x10 x10 1
               when x"00000034"   => data <= "11111110101101010001111011100011"; --bne x10 x11 -4
               when x"00000038"   => data <= "11111110101101010100100011100011"; --blt x10 x11 -16
               when x"0000003C"   => data <= "00000000011100000000000110010011"; --addi x3, x0 7
				-----------------------------------------------------------------------------------------
				------------------------------------------------------------------------------------------
				   --when x"00000000"   => data <= "00000000000000000000000100010011"; --addi x2 x0 0
               --when x"00000004"   => data <= "00000000000000010010010100000011"; --lw x10 0(x2)
               --when x"00000008"   => data <= "01000000000000000000010110010011"; --addi x11 x0 1024
               --when x"0000000C"   => data <= "00000000101001011100011000110011"; --xor x12,x11,x10
               --when x"00000010"   => data <= "11111110110001010000101011100011"; --beq x10,x12 loop
               --when x"00000014"   => data <= "11111110110001010000101011100011"; --beq x10,x12 loop
					--when x"00000018"   => data <= "01000000000000000000010110010011"; --addi x11 x0 1024
               --when x"0000001C"   => data <= "11111110010000010000000100010011"; --
               --when x"00000020"   => data <= "00000000101000010010011000100011"; --sw x10 12(x2)
               --when x"00000024"   => data <= "00000000110000010010011000000011"; --lw x12 12(x2)
               --when x"00000028"   => data <= "00000000000000000000010100010011"; --addi x10 x0 0
               --when x"0000002C"   => data <= "00000000101000000000010110010011"; --addi x11 x0 10
               --when x"00000030"   => data <= "00000000000101010000010100010011"; --addi x10 x10 1
               --when x"00000034"   => data <= "11111110101101010001111011100011"; --bne x10 x11 -4
               --when x"00000038"   => data <= "11111110101101010100100011100011"; --blt x10 x11 -16
               --when x"0000003C"   => data <= "00000000011100000000000110010011"; --addi x3, x0 7
					when x"00000040"   => data <= "00000000001000000000001000010011"; --addi x4,x0,2
					when x"00000044"   => data <= "00000000001100100111001100110011"; --and x6,x4,x3
					when x"00000048"   => data <= x"00000090";
					when x"0000004C"   => data <= x"00000090";
					when x"00000050"   => data <= x"00000090";
					when x"00000054"   => data <= x"00000090";
					when x"00000058"   => data <= x"00000090";
					when x"0000005C"   => data <= x"00000090";
					when x"00000060"   => data <= x"00000090";
					when x"00000064"   => data <= x"00000090";
					when x"00000068"   => data <= x"00000090";
					when x"0000006C"   => data <= x"00000090";
					when x"00000070"   => data <= x"00000090";
					when x"00000074"   => data <= x"00000090";
					when x"00000078"   => data <= x"00000090";
					when x"0000007C"   => data <= x"00000090";
					when x"00000080"   => data <= x"00000090";
               when others => data <= x"00000000";
            end case;
        end if;
    end process;
    

end architecture;